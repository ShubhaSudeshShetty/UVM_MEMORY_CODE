
package mem_pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "mem_sequence_item.sv"
`include "mem_sequence.sv"
`include "mem_sequencer.sv"
`include "mem_driver.sv"
`include "mem_monitor.sv"
`include "mem_agent.sv"
`include "mem_scoreboard.sv"
`include "mem_environment.sv"
`include "mem_test.sv"
endpackage
